library IEEE;
use IEEE.std_logic_1164.all;

package tankparameters is

constant  bullet_speed : integer := 5;
constant tank_height : integer := 30;
constant tank_width : integer := 60;
constant bullet_height : integer := 5;
constant bullet_width : integer := 5;

end package;



package body tankparameters is

end package body;
